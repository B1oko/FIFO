task clear;
    